module top(
    input clk
)


doublesha DUT


endmodule