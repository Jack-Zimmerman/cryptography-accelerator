module top(
    input logic CLK_100MHZ,
    input logic UART_TXD,
    output logic UART_RXD
);


//GLOBAL VARIABLES
logic rst_i; //global reset

//UART VARIABLES
logic finished_recieving; //status bit from UART rx
logic finished_sending; //status bit from UART tx
logic finished_read_byte; //byte completion for rx
logic finished_write_byte; //byte completion for tx
logic write_enable; //enable for UART tx
logic read_enable;
logic [7:0] read_bytes_passed; //we need to tally 608/8 = 76 bytes to read block info
logic [2:0] write_bytes_passed; //we need to tally 32/8 = 4 bytes to transmit nonce
logic [7:0] tx_byte; //feed buffer for tx
logic [7:0] rx_byte; //reciever buffer from rx
logic sending; //sending status bit

//TIMER VARIABLES
logic second_tick; //goes high when second has passed


//MINING VARIABLES
logic hash_enable; //enable for hashing 
logic [607:0] block_info; //everything needed for hashing besides nonce
logic [255:0] best_hash; //lowest hash achieved
logic [31:0] best_hash_nonce; //nonce corrosponding with best_hash




timer TIMER (
    .clk(CLK_100MHZ),
    .enable(hash_enable),
    .rst_i(rst_i),
    .second_tick(second_tick)
);

fsm FSM (
    .clk(CLK_100MHZ),
    .finished_recieving(finished_recieving),
    .finished_sending(finished_sending),
    .second_tick(second_tick),
    .rst_i(rst_i),
    .hash_enable(hash_enable),
    .write_enable(write_enable),
    .read_enable(read_enable)
);


hashcore HASHCORE (
    .clk(CLK_100MHZ),
    .enable(hash_enable),
    .rst_i(rst_i),
    .block_without_nonce(block_info),
    .best_hash(best_hash),
    .best_hash_nonce(best_hash_nonce)
);

uart_rx UART_RX(
    .i_Clock(CLK_100MHZ),
    .i_Rx_Serial(UART_RXD),
    .o_Rx_DV(finished_read_byte),
    .o_Rx_Byte(rx_byte)
);

uart_tx UART_TX (
    .i_Clock(CLK_100MHZ),
    .i_Tx_DV(write_enable),
    .i_Tx_Byte(tx_byte),
    .o_Tx_Active(sending),
    .o_Tx_Serial(UART_TXD),
    .o_Tx_Done(finished_write_byte)
);


always @(posedge CLK_100MHZ) begin
    //handle rx_byte
    if (read_enable) begin 
        if (finished_read_byte) begin
            if (read_bytes_passed == 8'd76) begin // we read the whole byte
                finished_recieving = 1; //set finish correctly
                read_bytes_passed = 0; 
            end else begin //otherwise read byte
                read_bytes_passed += 1;

                //serially load in block
                block_info[7:0] = rx_byte;
                block_info = block_info << 8;
            end
        end
    end else if (write_enable) begin
        if (finished_write_byte || write_bytes_passed == 3'b0) begin // we write the next byte
            if (write_bytes_passed == 3'd4) begin
                finished_sending = 1;
                write_bytes_passed = 0;
            end else begin //serially feed through the nonce
                tx_byte = best_hash_nonce[7:0];
                best_hash_nonce = best_hash_nonce << 8;

                write_bytes_passed += 1;
            end
        end 
    end
end


endmodule