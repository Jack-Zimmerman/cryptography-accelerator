module top(
    input logic CLK_100MHZ,
    input logic UART_TXD,
    output logic UART_RXD
);


fsm FSM (
    .
);


endmodule